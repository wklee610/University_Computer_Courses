`timescale 1ns/1ps

// 16에서 32비트로 변환
module signExtend(input[15:0] imm       
                , output[31:0] sign);       
    reg[31:0] trigger;          

    always @(imm) // input changes
        begin
            trigger <= 32'b1111_1111_1111_1111_0000_0000_0000_0000 + imm;           

            if(imm[15] == 0)            
            trigger <= 32'b0000_0000_0000_0000_0000_0000_0000_0000 + imm;           
        end
    assign sign = trigger; ////////////////// sign extension
endmodule

//////////////////// multi_plexers////////////////////
module big_mux(input wire[31:0] a                   
             , input wire[31:0] b               
             , input wire change                
             , output wire[31:0] result);               
    reg[31:0] trigger;

    always @({change,a,b}) ////////////////// change input
        begin
            trigger <= a;   

            if(change == 1) 
                trigger <= b;               
        end
    assign result = trigger;            
endmodule

module small_mux(input wire[4:0] a              
               , input wire[4:0] b              
               , input wire change                          
               , output wire[4:0] result);                  
    reg[4:0] trigger;           

    always @({change,a,b}) ////////////////// change input
        begin
            trigger <= a;

            if(change == 1)
                trigger <= b;
        end
    assign result = trigger;
endmodule

/////////////////////////////////// memory ///////////////////////////////////////
module MainMemory
    ( 
      input  CLOCK // clock
    , input  RESET // reset
    , input  ENABLE
    , input[31:0] FETCH_ADDRESS
    , input[64:0] EDIT_SERIAL

      //............../////////// Output
    , output reg[31:0] DATA
    );
  // /home/jimmy/VNMCC/src/MIPS/RAM.hs:40:1-7
  wire signed[63:0] c$wild_app_arg;
  wire  c$app_arg;
  // /home/jimmy/VNMCC/src/MIPS/RAM.hs:40:1-7
  wire signed[63:0] c$wild_app_arg_0;
  // /home/jimmy/VNMCC/src/MIPS/RAM.hs:40:1-7
  wire[63:0] a1;
  // /home/jimmy/VNMCC/src/MIPS/RAM.hs:40:1-7
  wire signed[63:0] wild;
  // /home/jimmy/VNMCC/src/MIPS/RAM.hs:40:1-7
  wire signed[63:0] wild_0;
  // /home/jimmy/VNMCC/src/MIPS/RAM.hs:40:1-7
  wire[63:0] ds;
  wire[31:0] c$i;

  assign c$wild_app_arg = $unsigned({{(64-32) {1'b0}},FETCH_ADDRESS});

  assign c$app_arg = EDIT_SERIAL[64:64] ? 1'b1 : 1'b0;

  assign c$i = ds[63:32];

  assign c$wild_app_arg_0 = $unsigned({{(64-32) {1'b0}},c$i});

  // blockRam begin
  reg[31:0] DATA_RAM[0:512-1];

  reg[16383:0] ram_init;
  integer i;
  initial begin
    ram_init = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
    for (i=0; i < 512; i = i + 1) begin
      DATA_RAM[512-1-i] = ram_init[i*32+:32];
    end
  end

  always @(posedge CLOCK) begin : DATA_blockRam

    if (c$app_arg & ENABLE) begin
      DATA_RAM[(wild_0)] <= ds[31:0]; //////////////////////
    end
    if (ENABLE) begin
      /////////////////////////////
      DATA <= DATA_RAM[(wild)]; /////////////
    end
  end
  // blockRam end 

  assign a1 = EDIT_SERIAL[63:0];

  assign wild = $signed(c$wild_app_arg);

  assign wild_0 = $signed(c$wild_app_arg_0);

  assign ds = EDIT_SERIAL[64:64] ? a1 : ({64 {1'bx}});


endmodule

/////////////////////////////// instruction ram ////////////////////////////////////
module InstructionRAM
    ( // Inputs
      input  CLOCK // clock
    , input  RESET // reset
    , input  ENABLE
    , input[31:0] FETCH_ADDRESS

      // Outputs
    , output reg[31:0] DATA
    );
  // /home/jimmy/VNMCC/src/MIPS/InstructionMem.hs:(17,1)-(23,30)
  wire signed[63:0] c$wild_app_arg;
  // /home/jimmy/VNMCC/src/MIPS/InstructionMem.hs:(17,1)-(23,30)
  wire signed[63:0] c$wild_app_arg_0;
  // /home/jimmy/VNMCC/src/MIPS/InstructionMem.hs:(17,1)-(23,30)
  wire[31:0] x1;
  // /home/jimmy/VNMCC/src/MIPS/InstructionMem.hs:(17,1)-(23,30)
  wire signed[63:0] wild;
  // /home/jimmy/VNMCC/src/MIPS/InstructionMem.hs:(17,1)-(23,30)
  wire signed[63:0] wild_0;
  wire[63:0] DATA_0;
  wire[63:0] x1_projection;

  assign c$wild_app_arg = $unsigned({{(64-32) {1'b0}},FETCH_ADDRESS});

  assign c$wild_app_arg_0 = $unsigned({{(64-32) {1'b0}},x1});

  assign DATA_0 = {64 {1'bx}};

  // blockRamFile begin
  reg[31:0] RAM[0:512-1];

  initial begin
    $readmemb("instructions.bin",RAM);
  end

  always @(posedge CLOCK) begin : InstructionRAM_blockRamFile
    if (1'b0 & ENABLE) begin
      RAM[(wild_0)] <= DATA_0[31:0];
    end
    if (ENABLE) begin
      DATA <= RAM[(wild)];
    end
  end
  // blockRamFile end

  assign x1_projection = {64 {1'bx}};

  assign x1 = x1_projection[63:32];

  assign wild = $signed(c$wild_app_arg);

  assign wild_0 = $signed(c$wild_app_arg_0);


endmodule

///////////////////////// ALU.v contents included below/////////////////////////
`include "ALU.v"



//iverilog -o out ALU.v

////////////// pipeline --> 5 stages total //////////////
module CPU(input wire RESET);
    integer i, j; // 

    wire[2:0] res_flags;
    wire[4:0] res_mux_rd;
    wire[31:0] res_inst
             , res_imm
             , res_mux_alu
             , res_alu
             , r_data
             , res_data_mem
             , res_brch
             , res_jmp;

    reg[31:0] register[31:0];
    reg[31:0] pc = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    reg CLOCK, ENABLE;

    reg ctrl_jmp = 0;
    
    reg[2:0] flags;
    //////////////////////////////// registers  
    reg[4:0] rs
           , rt
           , rd; 

    //////////////////////////////// opcode, function code  
    reg[5:0] opcode
           , func; 

    ///////////////////////////// main control
    reg[8:0] main_ctrl;
    
    
    reg[31:0] instruction
            , immediate;
    
    reg[31:0] reg_data_1
            , reg_data_2
            , w_data;

    //////////////////////////////// ALU    
    reg[31:0] alu_A
            , alu_B
            , mux_Alu_Out
            , Alu_Out;

    //////////////////////////////// pc  
    reg[31:0] pc_brch
            , pc_jmp
            , brch_Out
            , jmp_Out;

    //
    small_mux mux_readdata(rt
                         , rd
                         , main_ctrl[0]
                         , res_mux_rd);
    ////////////////////////////////
    big_mux mux_alu(reg_data_2
                  , immediate
                  , main_ctrl[1]
                  , res_mux_alu);

    big_mux mux_memory(Alu_Out
                     , r_data
                     , main_ctrl[7]
                     , res_data_mem);

    big_mux mux_branch(pc
                     , pc_brch
                     , {flags[0] & main_ctrl[5]}
                     , res_brch);

    big_mux mux_jump(brch_Out       
                     , pc_jmp                   
                     , ctrl_jmp         
                     , res_jmp);                


    signExtend mips_extend(instruction[15:0]
                         , res_imm);

    alu mips_alu(instruction
              , alu_A
              , alu_B
              , res_alu
              , res_flags);
    
    InstructionRAM mips_ram(CLOCK
                          , RESET
                          , ENABLE
                          , (pc)/4
                          , res_inst);
    
    MainMemory mips_memory(CLOCK
                         , RESET
                         , ENABLE
                         , {2'b00 , Alu_Out[31:2]}
                         , {main_ctrl[6], 2'b00 , Alu_Out[31:2] ,reg_data_2}
                         , r_data);



/////////////////////////////////////////////////////////////////////////////
    always @({RESET})
    begin
        for(i = 0; i < 99; i = i)
            begin
                CLOCK <= 1;                 
                ENABLE <= 1;                    
                register[0] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

                #10 //////////////////
                instruction <= res_inst;
                pc <= pc + 32'b0000_0000_0000_0000_0000_0000_0000_0100;

                #10 ////////////////// op_cd and func_cd
                opcode <= instruction[31:26];
                func <= instruction[5:0];

                    #10 //////////////////몰까
                    CLOCK <= 0;
                    
                    #10 //////////////////그로궤
                    CLOCK <= 1;

                #10 ////////////////// 메인 컨트롤
                if(opcode == 6'b000000 & func!=6'b001000)
                    begin
                        main_ctrl <= 10'b100001001; 
                        ctrl_jmp <= 0;
                    end
                /////////////////// R_instruction

                else if(opcode == 6'b001000 || opcode == 6'b001001 || opcode == 6'b001100 || opcode == 6'b001101 || opcode == 6'b001110 || opcode == 6'b001010 || opcode == 6'b001011 || opcode == 6'b001111) 
                    begin
                        main_ctrl <= 10'b100000010; 
                        ctrl_jmp <= 0;
                    end
                //////////////////// I_instruction

                else if(opcode == 6'b000010 || opcode == 6'b000011 || {opcode,func} == 12'b000000_001000)
                    begin
                        if(opcode == 6'b000011)
                            begin
                                register[31] <= pc;
                            end

                        pc_jmp <= {instruction[25:0],2'b00};
                        main_ctrl = 10'b000000000;
                        ctrl_jmp <= 1;
                    end
                //////////////////// J_instruction

                else if(opcode  ==  6'b000100  ||  opcode  ==  6'b000001 || opcode == 6'b000111 || opcode == 6'b000110 || opcode == 6'b000001 || opcode == 6'b000101)
                    begin
                        main_ctrl = 10'b000100100; 
                        ctrl_jmp <= 0;
                    end
                /////////////////// branch

                else if(opcode  ==  6'b100011 || opcode   ==   6'b100101 || opcode  ==  6'b100001 || opcode  ==  6'b100100 || opcode  ==  6'b100000 || opcode  ==  6'b100010 || opcode  ==  6'b100110)
                    begin
                        main_ctrl = 10'b110000010; 
                        ctrl_jmp <= 0;
                    end 
                ///////////////// 로드

                else if(opcode  ==  6'b101011 || opcode == 6'b101001 || opcode == 6'b101000 || opcode == 6'b101010 || opcode == 6'b101110)
                    begin
                        main_ctrl = 10'b001000010; 
                        ctrl_jmp <= 0;
                    end 
                ///////////////// 저장띠

                
                #10 ////////////// reg addr
                rs <= instruction[25:21];
                rt <= instruction[20:16];
                rd <= instruction[15:11];

                #10 //////////////// reg addr
                rd <= res_mux_rd;
                
                #10 ///////////////// reg Data
                reg_data_1 <= register[rs];
                reg_data_2 <= register[rt];

                    #10
                    CLOCK <= 0;
                    
                    #10
                    CLOCK <= 1;

                #10 /////////////// ALU Input
                alu_A <= reg_data_1;
                alu_B <= res_mux_alu;

                #10 /////////////// Jump reg
                if({opcode,func}  ==  12'b000000_001000)
                    pc_jmp <=  reg_data_1;

                #10 /////////////// ALU Output
                Alu_Out <= res_alu;
                flags <= res_flags;

                #10 /////////////// 16bit Immediate
                immediate <= res_imm;
                
                #10 /////////////// branch addr
                pc_brch <= pc + immediate<<2;

                    #10
                    CLOCK <= 0;
                    
                    #10
                    CLOCK <= 1;

                #10 ///////////////// write 2 memory
                if(main_ctrl[8]  ==  1'b1)
                    register[rd] <= res_data_mem;

                #10 ///////////////// branch
                brch_Out <= res_brch;
                CLOCK<=0;

                #10 ///////////////// jump
                pc <= res_jmp;
                ctrl_jmp <= 0;

                    #10
                    CLOCK <= 0;
                    
                    #10
                    CLOCK <= 1;

                #10 ///////////////// cpu end
                if(res_inst  ==  32'b1111_1111_1111_1111_1111_1111_1111_1111)
                    i = 99999999;
            end
            
            
            /////////////////////////// Display ///////////////////////////////
            for(j = 0; j < 512; j = j + 1)
                $display("%b", mips_memory.DATA_RAM[j]);
    end
endmodule