`timescale 1ns/1ps

module alu_test;

reg[31:0] Input, regA, regB;
wire[31:0] result;
wire[2:0] flags;


alu testalu(Input, regA, regB, result, flags);

initial begin
$display("Instructions RegA     RegB     Output   Flags");
$monitor("%h     %h %h %h %h %h %h",
Input, regA, regB, testalu.result, flags[0], flags[1], flags[2]);

    #10 
    //testing add 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1001;
    Input = 32'b000000_00000_00001_00000_00000_100000;


    #10 
    //testing addu 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_1111;
    Input = 32'b000000_00000_00001_00000_00000_100001;

    #10 
    //testing sub 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_1001;
    Input = 32'b000000_00000_00001_00000_00000_100010;

    #10 
    //testing subu 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB = 32'b0000_0000_0000_0000_0000_0000_1111_1111;
    Input = 32'b000000_00000_00001_00000_00000_100011;

    #10
    //testing and 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Input = 32'b000000_00000_00001_00000_00000_100100;

    #10
    //testing nor 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Input = 32'b000000_00000_00001_00000_00000_100111;

    #10
    //testing or 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Input = 32'b000000_00000_00001_00000_00000_100101;

    #10
    //testing xor 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
    Input = 32'b000000_00000_00001_00000_00000_100110;

    #10
    //testing addi 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1001;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b001000_00000_00001_0000000000000110;

    #10
    //testing addiu 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1001;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b001001_00000_00001_0000000000000110;

    #10
    //testing andi 
    regA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b001100_00000_00001_1111111111111111;

    #10
    //testing ori 
    regA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b001101_00000_00001_1111111111111111;

    #10
    //testing xori 
    regA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b100110_00000_00001_0000111100001111;

    #10
    //testing slt 
    regA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b000000_00000_00001_00000_00000_101010;

    #10
    //testing sltu 
    regA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b000000_00000_00001_00000_00000_101011;

    #10
    //testing slti 
    regA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b001010_00000_00001_0000000000001100;

    #10
    //testing sltiu 
    regA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b001011_00000_00001_0000000000001100;

    #10
    //testing sll 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    Input = 32'b000000_00000_00001_00000_01100_000000;

    #10
    //testing sllv 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    Input = 32'b000000_00000_00001_00000_01100_000100;

    #10
    //testing srl 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    Input = 32'b000000_00000_00001_00000_01100_000010;

    #10
    //testing srlv 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    Input = 32'b000000_00000_00001_00000_01100_000110;

    #10
    //testing sra 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    Input = 32'b000000_00000_00001_00000_01100_000011;

    #10
    //testing srav 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
    Input = 32'b000000_00000_00001_00000_01100_000111;

    #10
    //testing beq 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b000100_00000_00001_1111111111111111;

    #10
    //testing bne 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    Input = 32'b000101_00000_00001_1111111111111111;

    #10
    //testing lw 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1001;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    Input = 32'b100011_00000_00001_1111111111111111;

    #10
    //testing sw 
    regA = 32'b0000_0000_0000_0000_0000_0000_0000_1001;
    regB = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    Input = 32'b101011_00000_00001_1111111111111111;

#10 

$finish;

end

endmodule
